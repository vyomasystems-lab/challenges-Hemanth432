// See LICENSE.vyoma for details
module ALU_buggy(
  input [3:0]s,
  input ci, M,
  input [3:0] a, b,
  output reg [3:0] y
);

    reg [3:0] p, g;

    always @(*) begin

    p[0] <= ~(a[0] | (s[0] & b[0]) | (s[1] & ~b[0]));
    p[1] <= ~(a[1] | (s[0] & b[1]) | (s[1] & ~b[1]));
    p[2] <= ~(a[2] | (s[0] & b[3]) | (s[1] & ~b[2]));
    p[3] <= ~(a[3] | (s[0] & b[3]) | (s[1] & ~b[3]));

    g[0] <= ~((a[0] & ~b[0] & s[2]) | (a[0] & b[0] & s[3]));
    g[1] <= ~((a[1] & ~b[1] & s[2]) | (a[1] & b[1] & s[3]));
    g[2] <= ~((a[2] & ~b[2] & s[2]) | (a[2] & b[2] & s[3]));
    g[3] <= ~((a[3] & ~b[3] & s[2]) | (a[3] & b[3] & s[3]));

    y[0] = (p[0] ^ g[0]) ^ ~(~ci & ~M);
    y[1] = (p[1] ^ g[1]) ^ ~((~ci & ~M & g[0]) | (~M & p[0]));
    y[2] = (p[2] ^ g[2]) ^ ~((~ci & ~M & g[0] & g[1]) | (~M & p[1]) | (~M & p[0] & g[1]));
    y[3] = (p[3] ^ g[3]) ^ ~((~ci & ~M & g[0] & g[1] & g[2]) | (~M & p[2]) | (~M & p[1] & g[2]) | (~M & p[0] & g[1] & g[2]));
    end
endmodule